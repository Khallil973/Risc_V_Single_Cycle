module Alu_decoder (func3, func7, ALUOp,ALUControl,op5);
    input [6:0] op5, func7;
    input [2:0] func3;
    input [1:0] ALUOp;
    output [2:0] ALUControl;

    //interim wire
    wire [1:0] concatenation;

    assign concatenation = {op5[5], func7[5]};
    
    assign ALUControl = (ALUOp == 2'b00) ? 3'b000 :
                        (ALUOp == 2'b01) ? 3'b001 :
                        ((ALUOp == 2'b10) & (func3 == 3'b010)) ? 3'b101 :
                        ((ALUOp == 2'b10) & (func3 == 3'b110)) ? 3'b011 :
                        ((ALUOp == 2'b10) & (func3 == 3'b111)) ? 3'b010 :
                        ((ALUOp == 2'b10) & (func3 == 3'b000) & (concatenation == 2'b11)) ? 3'b001 :
                        ((ALUOp == 2'b10) & (func3 == 3'b000) & (concatenation != 2'b11)) ? 3'b000: 3'b000;

                        //We use != for rest of the 2bit condition like 00,01,10,and skip 11 condition
endmodule